--------------------------------------------------------------------------------
-- sw_interrupts.vhd: Demonstration of software interrupts implemented in
--                    hardware. Toggling of LEDs is generated via pressdown
--                    of buttons.
--
--                    Generics:
--                       - NUM_INTERRUPTS: The number of interrupt sources
--                                         (the number of buttons and LEDs).
--                    Inputs:
--                       - clock   : 50 MHz system clock.
--                       - reset_n : Inverting reset signal.
--                       - button_n: Push buttons for toggling leds.
--                    Outputs:
--                       - led     : LEDs toggled by pressdown of the buttons.
--
--                    Hardware implemented for FPGA card Terasic DE0.
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sw_interrupts is
   generic(NUM_INTERRUPTS: natural range 1 to 3 := 3);
   port(clock, reset_n   : in std_logic;
        button_n         : in std_logic_vector(NUM_INTERRUPTS - 1 downto 0); 
        led              : out std_logic_vector(NUM_INTERRUPTS - 1 downto 0));
end entity;

architecture behaviour of sw_interrupts is
signal led_s: std_logic_vector(NUM_INTERRUPTS - 1 downto 0);
begin

   --------------------------------------------------------------------------------
   -- OUTPUT_PROCESS: Toggling LEDs at pressdown of corresponding push buttons.
   --                 Edge detection is generated by comparing current input
   --                 signals with previous input signals, stored via a variable.
   --                 This happens at rising edge of the clock. All LEDs are
   --                 disabled at system reset.
   --------------------------------------------------------------------------------
   OUTPUT_PROCESS: process(clock, reset_n) is
   variable button_previous_n: std_logic_vector(NUM_INTERRUPTS - 1 downto 0);
   begin
      if (reset_n = '0') then
         led_s <= (others => '0');
         button_previous_n := (others => '1');
      elsif (rising_edge(clock)) then
         for i in 0 to NUM_INTERRUPTS - 1 loop
            if (button_n(i) = '0' and button_previous_n(i) = '1') then
               led_s(i) <= not led_s(i);
            end if;
         end loop;
      button_previous_n := button_n;
      end if;
   end process;
   
   led <= led_s;

end architecture;